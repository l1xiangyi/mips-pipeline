`include "alu.v"
`timescale 1ns/1ps

module alu_test;

reg[31:0] instruction,regA,regB;
wire[31:0] result;
wire[2:0] flags;

alu testalu(instruction, regA, regB, result, flags);

task test_bench;
    input[31:0] instruction_t;
    input[31:0] regA_t, regB_t;
    input[31:0] result_t;
    input[2:0] flags_t;
    begin
        instruction = instruction_t;
        regA = regA_t;
        regB = regB_t;
        #10
        $write("instruction:%b; regA:%h regB:%h opcode:%h funct:%h; result:%h flags:%b;\tInfo: ",instruction_t,regA_t,regB_t,testalu.opcode,testalu.funct,result,flags);
        if(result === result_t && flags === flags_t)
            $display("PASS");
        else
            $display("WRONG");       
    end
endtask

initial begin

#10 $display("add");
#10 test_bench(32'b000000_00001_00000_00000_00000_100000,-2,2,8'b00000000,3'b100); // -2+2=0
#10 test_bench(32'b000000_00001_00000_00000_00000_100000,32'h80000001,32'h80000001,32'h00000002,3'b001); //10...01+10...01=0...10 overflow
#10 test_bench(32'b000000_00001_00000_00000_00000_100000,32'h7ffffffe,32'h00000002,32'h80000000,3'b001); // 01...10+0...010=10...0 overflow

#10 $display("\naddi");
#10 test_bench(32'b001000_00000_00001_1111111111111110,3,32'bx,1,3'b000);//-2+3=1
#10 test_bench(32'b001000_00000_00001_1000000000000000,32'h80000000,32'bx,32'h7fff8000,3'b001);//10...0+1...10...0=01...10...0 overflow
#10 test_bench(32'b001000_00000_00001_0000000000000010,32'h7ffffffe,32'bx,32'h80000000,3'b001); //01...10+0...010=10...0 overflow 
#10 test_bench(32'b001000_00000_00001_0000000000000010,-3,32'bx,-1,3'b000);

#10 $display("\naddu");
#10 test_bench(32'b000000_00001_00000_00000_00000_100001,-2,2,0,3'b100);
#10 test_bench(32'b000000_00001_00000_00000_00000_100001,-2147483647,-2147483647,2,3'b000);
#10 test_bench(32'b000000_00001_00000_00000_00000_100001,2147483647,1,32'h80000000,3'b000);
#10 test_bench(32'b000000_00001_00000_00000_00000_100001,7,8,15,3'b000);

#10 $display("\naddiu");
#10 test_bench(32'b001001_00000_00001_0000000000000111,8,32'bx,15,3'b000);
#10 test_bench(32'b001001_00000_00001_1000000000000000,32'h80000000,32'bx,32'h7fff8000,3'b000);


#10 $display("\nsub");
#10 test_bench(32'b000000_00001_00000_00000_00000_100010,2,-2,4,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00000_100010,-2147483647,2,32'h7fffffff,3'b001);
#10 test_bench(32'b000000_00000_00001_00000_00000_100010,32'h7fffffff,-1,32'h80000000,3'b001);


#10 $display("\nsubu");
#10 test_bench(32'b000000_00000_00001_00000_00000_100011,-2147483647,2,32'h7fffffff,3'b000);
#10 test_bench(32'b000000_00001_00000_00000_00000_100011,2147483646,-2,32'h8000_0000,3'b000);

#10 $display("\nand");
#10 test_bench(32'b000000_00001_00000_00000_00000_100100,32'h00000001,32'h11111111,32'h0000_0001,3'b000);

#10 $display("\nandi");
#10 test_bench(32'b001100_00000_00001_0000000000000001,32'hffffffff,32'bx,32'h00000001,3'b000);

#10 $display("\nnor");
#10 test_bench(32'b000000_00001_00000_00000_00000_100111,32'h00000001,32'h00000010,32'hffffffee,3'b000);

#10 $display("\nori");
#10 test_bench(32'b001101_00000_00001_0000000000000001,32'h00000010,32'bx,32'h00000011,3'b000);

#10 $display("\nxor");
#10 test_bench(32'b000000_00001_00000_00000_00000_100110,32'b00000001,32'b00000011,32'b00000010,3'b000);

#10 $display("\nxori");
#10 test_bench(32'b001110_00000_00001_0000000000000001,32'b00000011,32'bx,32'b00000010,3'b000);

#10 $display("\nbeq");
#10 test_bench(32'b000100_00001_00000_1000000000100000,2,2,32'b0,3'b100);
#10 test_bench(32'b000100_00000_00001_1000000000100000,3,2,32'b1,3'b000);

#10 $display("\nbne");
#10 test_bench(32'b000101_00001_00000_1000000000100000,2,2,32'b0,3'b100);
#10 test_bench(32'b000101_00000_00001_1000000000100000,3,2,32'b1,3'b000);

#10 $display("\nslt");
#10 test_bench(32'b000000_00000_00001_00000_00000_101010,-5,-1,32'h00000001,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00000_101010,5,5,32'h00000000,3'b100);
#10 test_bench(32'b000000_00000_00001_00000_00000_101010,8,-9,32'h00000001,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00000_101010,-9,8,32'h00000000,3'b100);

#10 $display("\nslti");
#10 test_bench(32'b001010_00000_00001_1000000000000001,2,2,0,3'b100); // 1000000000000001 = -32767
#10 test_bench(32'b001010_00000_00001_0000000000000101,3,3,1,3'b000);
#10 test_bench(32'b001010_00000_00001_1111111111111111,-3,-3,1,3'b000);
#10 test_bench(32'b001010_00000_00001_0111111111111111,-3,-3,1,3'b000);

#10 $display("\nsltiu");
#10 test_bench(32'b001011_00000_00001_1111111111111111,3,3,1,3'b000); // 1111111111111111 = -1
#10 test_bench(32'b001011_00000_00001_0111111111111111,-3,-3,0,3'b100); // -3 = 1111111111111101

#10 $display("\nsltu");
#10 test_bench(32'b000000_00001_00000_00000_00000_101011,-1,-3,0,3'b100); 
#10 test_bench(32'b000000_00001_00000_00000_00000_101011,-3,-1,1,3'b000);

#10 $display("\nlw");
#10 test_bench(32'b100011_00001_00000_1111111111111111,32'bx,-3,-4,3'b000);
#10 test_bench(32'b100011_00001_00000_0000000000000011,32'bx,2,5,3'b000);

#10 $display("\nsw");
#10 test_bench(32'b101011_00001_00000_1111111111111111,32'bx,-3,-4,3'b000);
#10 test_bench(32'b101011_00001_00000_0000000000000011,32'bx,2,5,3'b000);

#10 $display("\nsll");
#10 test_bench(32'b000000_00001_00000_00000_00010_000000,1,1,4,3'b000);
#10 test_bench(32'b000000_00001_00000_00000_00011_000000,32'h111,32'h111,32'h888,3'b000);

#10 $display("\nsllv");
#10 test_bench(32'b000000_00000_00001_00000_00000_000100,4,1,16,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00000_000100,4,3,48,3'b000);

#10 $display("\nsrl");
#10 test_bench(32'b000000_00000_00001_00000_00010_000010,32'bx,8,2,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00011_000010,32'bx,2,0,3'b100);

#10 $display("\nsrlv");
#10 test_bench(32'b000000_00000_00001_00000_00000_000110,2,8,2,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00000_000110,3,15,1,3'b000);

#10 $display("\nsra");
#10 test_bench(32'b000000_00000_00001_00000_00010_000011,32'bx,8,2,3'b000);
#10 test_bench(32'b000000_00000_00001_00000_00100_000011,32'bx,32'hffffff00,32'hfffffff0,3'b000);

#10 $display("\nsrav");
#10 test_bench(32'b000000_00000_00001_00000_00000_000111,4,32'hf,0,3'b100);
#10 test_bench(32'b000000_00000_00001_00000_00000_000111,4,32'h80000000,32'hf8000000,3'b000);


#10 $finish;

end

endmodule