// CLK: input clock signal

module CPU
(
    //input
      input CLK
);